module init_values_loader (
    clk, rst, center_peek, l, w
)
input

endmodule