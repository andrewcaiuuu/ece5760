module single_node_zero_inital(

);

endmodule