

module xy2addr(

)

endmodule