module init_values_LUT (
    output reg [17:0] node_value_out,
    input wire [18:0] address
);

reg [17:0] node_values [0:29];

initial
begin
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0C924
    0x0DB6D
    0x0DB6D
    0x0DB6D
    0x0DB6D
    0x0DB6D
    0x0DB6D
    0x0C924
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0C924
    0x0DB6D
    0x0EDB6
    0x0EDB6
    0x0EDB6
    0x0EDB6
    0x0DB6D
    0x0C924
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0C924
    0x0DB6D
    0x0EDB6
    0x10000
    0x10000
    0x0EDB6
    0x0DB6D
    0x0C924
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0C924
    0x0DB6D
    0x0EDB6
    0x10000
    0x10000
    0x0EDB6
    0x0DB6D
    0x0C924
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0C924
    0x0DB6D
    0x0EDB6
    0x0EDB6
    0x0EDB6
    0x0EDB6
    0x0DB6D
    0x0C924
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0C924
    0x0DB6D
    0x0DB6D
    0x0DB6D
    0x0DB6D
    0x0DB6D
    0x0DB6D
    0x0C924
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0C924
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0B6DB
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x0A492
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x09249
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x08000
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x06DB6
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x05B6D
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x04924
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x036DB
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x02492
    0x01249
    0x00000
    0x00000
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x01249
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000
    0x00000

end

always @(address)
begin
    if (address < 30)
        node_value_out = node_values[address];
    else
        node_value_out = 18'h00000;
end

endmodule