module solver()